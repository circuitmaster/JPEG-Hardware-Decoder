//////////////////////////////////////////////////////////////////////////////////
// Module Name: Number Generator
// Description: Generates number from endecoded image sequence
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module Number_Generator(
    input clk, rst
);
    
    
    
endmodule